// Matrix Multiplication Accelerator
`timescale 1ns / 1ps

module matrix_mul (
    input wire clk,
    input wire rst_n,
    input wire [7:0] matrix_a [15:0],
    input wire [7:0] matrix_b [15:0],
    input wire start,
    output reg done,
    output reg [15:0] result [15:0]
);

    // State machine
    localparam IDLE = 2'b00;
    localparam COMPUTE = 2'b01;
    localparam DONE = 2'b10;

    reg [1:0] state;
    reg [3:0] i, j, k;
    reg [15:0] temp_result;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            done <= 1'b0;
            i <= 4'b0;
            j <= 4'b0;
            k <= 4'b0;
        end else begin
            case (state)
                IDLE: begin
                    if (start) begin
                        state <= COMPUTE;
                        i <= 4'b0;
                        j <= 4'b0;
                        k <= 4'b0;
                    end
                end

                COMPUTE: begin
                    if (i < 4) begin
                        if (j < 4) begin
                            if (k < 4) begin
                                temp_result <= temp_result + 
                                    matrix_a[i*4 + k] * matrix_b[k*4 + j];
                                k <= k + 1;
                            end else begin
                                result[i*4 + j] <= temp_result;
                                temp_result <= 16'b0;
                                k <= 4'b0;
                                j <= j + 1;
                            end
                        end else begin
                            j <= 4'b0;
                            i <= i + 1;
                        end
                    end else begin
                        state <= DONE;
                        done <= 1'b1;
                    end
                end

                DONE: begin
                    if (!start) begin
                        state <= IDLE;
                        done <= 1'b0;
                    end
                end
            endcase
        end
    end

endmodule
